`default_nettype none

// just a stub to keep the Tiny Tapeout tools happy

module tt_um_tkmdemo (
    input  wire       VGND,
    input  wire       VPWR,
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    inout  wire [7:0] ua, // analog pins
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);
    assign uio_out = 0;
    assign uio_oe = 0;
    assign uo_out(0) = ui_in[0] ^ ui_in[1]; 
    assign uo_out(0) = ui_in[0] & ui_in[1];
    assign uo_out[7:2] =6'b0;
    
    
    
    

endmodule
